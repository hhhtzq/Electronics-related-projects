    Mac OS X            	   2  �     �                                    ATTR;���  �  $   �                 $     com.apple.TextEncoding     3     com.apple.lastuseddate#PS      C   H  com.apple.macl #   �   Y  7com.apple.metadata:kMDLabel_7e3pzpa3rf3xsfxrvvtgdhvs6i  utf-8;134217984���^    Gu5#     �:��=G������H� �޲�F���V���                                    �$�c�m[[p�6��vI�H�ҧkDp���4� ���ת7�}Y�j�9l�6�R��`�l�Wfa��Q��ȩ���g��kĸ�g�b4�K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           This resource fork intentionally left blank                                                                                                                                                                                                                            ��